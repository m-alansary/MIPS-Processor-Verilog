module register



endmodule
